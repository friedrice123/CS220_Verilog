always @(result) begin
    //     $display("result=%d",a);
    // end