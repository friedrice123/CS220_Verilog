module instruction_memory(address, instruction);
    input [31:0] address;
    output [31:0] instruction;

    reg [31:0] memory[0:15];

    initial begin
        memory[0]= 32'b000000_00000_00001_00010_00000_100000;
        memory[1]= 32'b000000_00000_00001_00011_00000_100011;
        memory[2]= 32'b000000_00000_00001_00100_00000_100100;
        memory[3]= 32'b000000_00000_00001_00101_00000_100101;
        memory[4]= 32'b000000_00000_00001_00110_00010_000000;
        memory[5]= 32'b000000_00000_00001_00110_00000_100101;
        memory[6]= 32'b000101_00000_00001_00000_00000_001000;
        memory[7]= 32'b010100_00000_00000_00000_00000_001000;
        memory[8]= 32'b001000_00000_00000_00000_00000_100000;
        memory[9]= 32'b000000_00000_00000_00000_00000_000000;
        memory[10]=32'b000000_00000_00000_00000_00000_000000;
        memory[11]=32'b000000_00000_00000_00000_00000_000000;
        memory[12]=32'b000000_00000_00000_00000_00000_000000;
        memory[13]=32'b000000_00000_00000_00000_00000_000000;
        memory[14]=32'b000000_00000_00000_00000_00000_000000;
        memory[15]=32'b000000_00000_00000_00000_00000_000000;
    end
    
    assign instruction=memory[address];
endmodule