`include "floating_point_addition.v" 
module test;
reg [31:0] a,b;
wire [31:0]sum;
floatAdder uut (.a(a),.b(b),.sum(sum));
initial begin
    a=32'b0_10000101_10100101110011001100110; //105.45
    b=32'b0_10000011_01100101000111101011100; //22.32
    #100;
    $display("%b",sum);//127.77
    #100;
    a=32'b0_10000101_10100101110011001100110; //105.45
    b=32'b1_10000011_01100101000111101011100; //-22.32
    #100;
    $display("%b",sum);//83.13
    a=32'b01000000101101010111000010100100; //5.67
    b=32'b11000001111001110000101000111101; //-28.88
    #100;
    $display("%b",sum);//-23.21
    a=32'b11000000101101010111000010100100; //-5.67
    b=32'b11000001111001110000101000111101; //-28.88
    #100;
    $display("%b",sum);//-34.55
    $finish;
end
endmodule