module something (
    
);
    
endmodule